///////////////////////////////////////////////////////////////////////////////////
// Testbench for Component: MUX4
// Package: FIUSCIS-CDA
// Course: CDA3102 (Computer Architecture), Florida International University
// Developer: Trevor Cickovski
// License: MIT, (C) 2020 All Rights Reserved
///////////////////////////////////////////////////////////////////////////////////


module testbench();
`include "../Test/Test.v"

///////////////////////////////////////////////////////////////////////////////////
// Inputs: A, B, C, D (1-bit), S (2-bit)
reg A, B, C, D;
reg[1:0] S;
///////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////
// Output: Y (1-bit)
wire Y;
///////////////////////////////////////////////////////////////////////////////////

MUX4 myMUX(A, B, C, D, S, Y);

initial begin
////////////////////////////////////////////////////////////////////////////////////////
// Test: S=00
$display("Testing: S=00");
A=1; B=0; C=0; D=0; S=2'b00;  #10; 
verifyEqual(Y, A);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: S=01
$display("Testing: S=01");
A=0; B=1; C=0; D=0; S=2'b01;  #10; 
verifyEqual(Y, B);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: S=10
$display("Testing: S=10");
A=0; B=0; C=1; D=0; S=2'b10;  #10; 
verifyEqual(Y, C);
////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////
// Test: S=11
$display("Testing: S=11");
A=0; B=0; C=0; D=1; S=2'b11;  #10; 
verifyEqual(Y, D);
////////////////////////////////////////////////////////////////////////////////////////
$display("All tests passed.");
end

endmodule